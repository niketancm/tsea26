
module adder_ctrl
  (
    input wire [2:0]    function_i,
    input wire 		opa_sign_i,
    output wire 	mx_opa_inv_o,
    output wire [1:0] 	mx_ci_o
   );

   // Remove the following lines and put your code here
   assign 		mx_opa_inv_o = 0;
   assign 		mx_ci_o = 0;

endmodule // adder_ctrl
