
module min_max_ctrl
  (
    input wire [2:0]    function_i,
    input wire 		opa_sign_i,
    input wire 		opb_sign_i,
    input wire 		carry_i,
    output wire 	mx_minmax_o
   );

   // Remove the following line and put your code here
   assign 		mx_minmax_o = 0;

endmodule // min_max_ctrl
